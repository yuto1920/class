module strange(
  input  wire       clk,
  input  wire       res,
  input  wire [1:0] s,
  output reg  [1:0] state
);

/* ���̕����ɁA�K�v�ȉ�H���������݂܂��傤 */

endmodule

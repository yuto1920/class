module mult2 (
  input  wire [3:0] a,
  input  wire [3:0] b,
  output wire [7:0] mult
);

/* ���̕����ɕK�v�ȉ�H���L�q���Ă��������B*/

endmodule
